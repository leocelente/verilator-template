module top;
/* 
  Module: Top
  Description: This is a test module to test a SystemVerilog Simulation
  toolchain based on Verilator
*/
initial begin 
  
  $display("\n\n\tHello World\n"); 
  $finish; 
  
end
endmodule
